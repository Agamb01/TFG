----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:22:59 01/07/2015 
-- Design Name: 
-- Module Name:    main - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity main is
end main;

architecture Behavioral of main is
----------------------------Instruction Fetch-----------------------------
----------------------------Instruction Fetch-----------------------------

----------------------------Instruction Decode----------------------------
----------------------------Instruction Decode----------------------------

---------------------------------Execution--------------------------------
---------------------------------Execution--------------------------------

----------------------------------Memory----------------------------------
----------------------------------Memory----------------------------------

--------------------------------Write Back--------------------------------
--------------------------------Write Back--------------------------------

begin

----------------------------Instruction Fetch-----------------------------
----------------------------Instruction Fetch-----------------------------

----------------------------Instruction Decode----------------------------
----------------------------Instruction Decode----------------------------

---------------------------------Execution--------------------------------
---------------------------------Execution--------------------------------

----------------------------------Memory----------------------------------
----------------------------------Memory----------------------------------

--------------------------------Write Back--------------------------------
--------------------------------Write Back--------------------------------


end Behavioral;

