----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:47:54 01/22/2015 
-- Design Name: 
-- Module Name:    EXE_main - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- Entradas:
--    Clock de sistema
--    Reset de sistema
--    Array de paradas de la siguiente instrucci�n
--    Bit de instruccion "NULA" siguiente

--    Contador de programa para calcular direccion de salto
--    Entero sacado de la instruccion
--    Buses de datos de los registros seleccionados por la instruccion

--    Se�ales de control para etapa de ejecucion:
--       bits[3:1] -> ALU_op
--       bits[0]   -> ALU_ctr

-- Salidas:
--    Array de paradas de esta instrucci�n
--    Bit de instrucci�n "NULA" actual
--    Enable para l�gica de fase

--    Direccion de salto calculada
--    Resultado de operacion calculado por la ALU
--    Flags de la operacion calculada por la ALU

library work;
   use work.my_package.all;
   
entity EXE_main is
   Port( 
      clk, rst       : in STD_LOGIC;
            
      --Entradas (ID->EXE)
      in_PC          : in STD_LOGIC_VECTOR(31 downto 0);
      in_entero      : in STD_LOGIC_VECTOR(31 downto 0);
      in_busA        : in STD_LOGIC_VECTOR(31 downto 0);
      in_busB        : in STD_LOGIC_VECTOR(31 downto 0);
       
      --Salidas (EXE->MEM)
      out_PC_salto   : out STD_LOGIC_VECTOR(31 downto 0);
      out_ALU_bus    : out STD_LOGIC_VECTOR(31 downto 0);
      out_ALU_flags  : out STD_LOGIC_VECTOR(1 downto 0); -- Flags(N,Z)

      --Se�ales de control(ID->EXE)
      in_EXE_control : in STD_LOGIC_VECTOR(3 downto 0);
        -- [3:1]=ALUop, [0]=ALUsrc

   -- Entradas y salidas de paso, sirven para simplificar el dise�o superior
      in_regW         : in STD_LOGIC_VECTOR(3 downto 0);  -- Registro destino
      in_WB_control   : in STD_LOGIC_VECTOR(1 downto 0);
      in_MEM_control  : in STD_LOGIC_VECTOR(5 downto 0);
      
      out_BusB        : out STD_LOGIC_VECTOR(31 downto 0);
      out_regW        : out STD_LOGIC_VECTOR(3 downto 0);  -- Registro destino
      out_WB_control  : out STD_LOGIC_VECTOR(1 downto 0);
      out_MEM_control : out STD_LOGIC_VECTOR(5 downto 0)

   );
end EXE_main;

architecture Behavioral of EXE_main is

-- Modulo que realiza el trabajo de la fase
   component Phase2_Execution is
      port (  
         --Entradas (ID->EXE)
         in_PC          : in STD_LOGIC_VECTOR(31 downto 0);
         in_entero      : in STD_LOGIC_VECTOR(31 downto 0);
         in_busA        : in STD_LOGIC_VECTOR(31 downto 0);
         in_busB        : in STD_LOGIC_VECTOR(31 downto 0);
          
         --Salidas (EXE->MEM)
         out_PC_salto   : out STD_LOGIC_VECTOR(31 downto 0);
         out_ALU_bus    : out STD_LOGIC_VECTOR(31 downto 0);
         out_ALU_flags  : out STD_LOGIC_VECTOR(1 downto 0); -- Flags(N,Z)

         --Se�ales de control(ID->EXE)
         in_EXE_control : in STD_LOGIC_VECTOR(3 downto 0) 
           -- [3:1]=ALUop, [0]=ALUsrc
      );
   end component;

   signal s_ALU_flags     : STD_LOGIC_VECTOR(1 downto 0); -- Flags(N,Z)
   signal s_ALU_flags_reg : STD_LOGIC_VECTOR(1 downto 0); -- Flags(N,Z)

begin

-- Se�ales de paso, sirven para simplificar el dise�o superior
   out_regW        <= in_regW;
   out_WB_control  <= in_WB_control;
   out_MEM_control <= in_MEM_control;
   out_BusB        <= in_BusB;
      
-- Modulo funcional de la fase EXE
   i_pEXE: Phase2_Execution
      Port map (
         --Entradas (ID->EXE)
         in_PC => in_PC,
         in_entero => in_entero,
         in_busA => in_busA,
         in_busB => in_busB,
         
         --Salidas (EXE->MEM)
         out_PC_salto => out_PC_salto,
         out_ALU_bus => out_ALU_bus,
         out_ALU_flags => s_ALU_flags,

         --Se�ales de control(ID->EXE)
         in_EXE_control => in_EXE_control
      );

--Registro flags
   out_ALU_flags <= s_ALU_flags_reg;

   --Proceso guarda flags en registros
   p_arith: process(clk, rst)
   begin
      if rst='0' then 
         s_ALU_flags_reg <= "00";
      elsif rising_edge(clk) then
         if in_EXE_control(3 downto 1) = "111" then
            s_ALU_flags_reg <= s_ALU_flags;
         end if;
      end if;
   end process;
   
end Behavioral;

